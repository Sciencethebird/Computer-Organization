//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:    0511105   
//----------------------------------------------
//Date:     2019/05/23
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
//reg     [32-1:0] data_o;

//Sign extended
assign data_o[31:16] = (data_i[15] == 0) ? 16'h0000 : 16'hffff;
assign data_o[15:0] = data_i[15:0];
          
endmodule      
     